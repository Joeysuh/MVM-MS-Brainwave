/***************************************************/
/* ECE 327: Digital Hardware Systems - Spring 2025 */
/* Lab 4                                           */
/* MVM Control FSM                                 */
/***************************************************/

module ctrl # (
    parameter VEC_ADDRW = 8,
    parameter MAT_ADDRW = 9,
    parameter VEC_SIZEW = VEC_ADDRW + 1,
    parameter MAT_SIZEW = MAT_ADDRW + 1
    
)(
    input  clk,
    input  rst,
    input  start,
    input  [VEC_ADDRW-1:0] vec_start_addr, // vector start addr
    input  [VEC_SIZEW-1:0] vec_num_words, // size of vec in word (4)
    input  [MAT_ADDRW-1:0] mat_start_addr, // matrix start addr
    input  [MAT_SIZEW-1:0] mat_num_rows_per_olane, // num of rows assigned to each olane.
    output [VEC_ADDRW-1:0] vec_raddr, // vector read addr - generated by controller
    output [MAT_ADDRW-1:0] mat_raddr, // matrix read addr - generated by controller
    output accum_first, // signals first compute
    output accum_last, // signals last compute
    output ovalid,
    output busy 
);

/******* Your code starts here *******/
enum {IDLE, COMPUTE} state, next_state;

logic [VEC_ADDRW-1:0] vec_start_addr_r; // wire for vec start
logic [VEC_SIZEW-1:0] vec_num_words_r; // vec word size
logic [MAT_ADDRW-1:0] mat_start_addr_r; // wire for mat start
logic [MAT_SIZEW-1:0] mat_num_rows_per_olane_r; // rows per olane

// Internal output wires
logic [VEC_ADDRW-1:0] vec_raddr_r;
logic [MAT_ADDRW-1:0] mat_raddr_r;
logic accum_first_r;
logic accum_last_r;
logic ovalid_r;
logic busy_r;

// reg for output addr
logic [VEC_ADDRW-1:0] vec_raddr_out_reg;
logic [MAT_ADDRW-1:0] mat_raddr_out_reg;

// counters to locate where we are
logic [VEC_SIZEW-1:0] word_counter;
logic [MAT_SIZEW-1:0] row_counter;

always_ff @(posedge clk) begin
    if (rst) begin
        state <= IDLE;
        vec_start_addr_r <= 0;
        vec_num_words_r <= 0;
        mat_start_addr_r <= 0;
        mat_num_rows_per_olane_r <= 0;
        word_counter <= 0;
        row_counter <= 0;

        // reset output registers
        vec_raddr_r <= 0;
        mat_raddr_r <= 0;
        accum_first_r <= 0;
        accum_last_r <= 0;
        ovalid_r <= 0;
        busy_r <= 0;

    end else begin
        state <= next_state;

        if (state == IDLE) begin
            if (start) begin
                vec_start_addr_r <= vec_start_addr;
                vec_num_words_r <= vec_num_words;
                mat_start_addr_r <= mat_start_addr;
                mat_num_rows_per_olane_r <= mat_num_rows_per_olane;
                word_counter <= 0;
                row_counter <= 0;
            end
            
            vec_raddr_r <= 0;
            mat_raddr_r <= 0;
            accum_first_r <= 0;
            accum_last_r <= 0;
            ovalid_r <= 0;
            busy_r <= 0;
        end else if (state == COMPUTE) begin
            vec_raddr_r <= vec_start_addr_r + word_counter;
            mat_raddr_r <= mat_start_addr_r + row_counter * vec_num_words_r + word_counter;
            ovalid_r <= 1;
            busy_r <= 1;
            if (word_counter == 0) begin
                accum_first_r <= 1;
            end else begin
                accum_first_r <= 0;
            end
            if (word_counter == vec_num_words_r - 1) begin
                accum_last_r <= 1;
            end else begin
                accum_last_r <= 0;
            end
            // counter 
            if (word_counter == vec_num_words_r - 1) begin
                word_counter <= 0;
                row_counter  <= row_counter + 1;
            end else begin
                word_counter <= word_counter + 1;
            end
        end
    end
end


always_comb begin: state_decoder
    case (state) 
        IDLE: begin
            if (start) next_state = COMPUTE; else next_state = IDLE;
        end
        
        COMPUTE: begin
            if ((word_counter == vec_num_words_r -1) && (row_counter == mat_num_rows_per_olane_r -1)) begin 
                next_state = IDLE;
            end else 
                next_state = COMPUTE;
        end
        default: next_state = IDLE;
    endcase
end


assign vec_raddr = vec_raddr_r;
assign mat_raddr = mat_raddr_r;
assign accum_first = accum_first_r;
assign accum_last = accum_last_r;
assign ovalid = ovalid_r;
assign busy = busy_r;


/******* Your code ends here ********/

endmodule